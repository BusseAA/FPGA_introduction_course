module counter #(
	parameter BW_VAL = 16,
	parameter MAX_VAL = 2
)(
	input clk,
	output [BW_VAL-1: 0] val
);

reg [BW_VAL-1: 0] cnt;

/*
*	counter code and input/output connection
*/

endmodule