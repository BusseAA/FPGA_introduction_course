module top(
	input CLK,
	output DS_EN1, DS_EN2, DS_EN3, DS_EN4,
	output DS_A, DS_B, DS_C, DS_D, DS_E, DS_F, DS_G
);

	wire [3:0] d = 4'b1010;
	wire [3:0] anodes;
	assign {DS_EN1, DS_EN2, DS_EN3, DS_EN4} = ~anodes;
	
	wire [6:0] segments;
	assign {DS_A, DS_B, DS_C, DS_D, DS_E, DS_F, DS_G} = segments; // for some boards you should invert segments (~segments)
	
	clk_div clk_div(.clk(CLK), .clk2(clk2));
	bin_display disp(.clk(clk2), .data(d), .anodes(anodes), .segments(segments));
	
endmodule